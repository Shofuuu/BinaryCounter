library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity BinaryCounter_top is
  Port (
    clk: in STD_LOGIC;
    led: out STD_LOGIC_VECTOR (7 to 0)
  );
end entity;

architecture BinaryCounter_top of BinaryCounter_top is
begin

end architecture;
